module main
import crayon

fn corpus() {

}

fn grineer() {
	
}